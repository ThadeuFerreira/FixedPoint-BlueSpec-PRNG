package InterfaceLogTableFxdP;

interface InterfaceLogTableFxdP#(
   type input_type,
   type out_type
);

   method out_type get (input_type i);
 
endinterface: InterfaceLogTableFxdP

endpackage: InterfaceLogTableFxdP